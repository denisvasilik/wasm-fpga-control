library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

package WasmFpgaControlPackage is

end package;

package body WasmFpgaControlPackage is

end package body;
